
module EX(
    input       clk,
    input       rst,

    input   [31:0] alu1_ex_in,
    input   [31:0] alu2_ex_in,
    input   [4:0]  ALUOp,

    input   [31:0] pc_ex_in,
    input   [31:0] imm_ex_in,
    input   [2:0] NPCOp_ex_in,

    input       MemWrite_ex_in,
    input       DMType_ex_in,
    input       
);

endmodule